
input [7:0] tmp;
input [3:0] cnt;

assign 

always @(*) begin
    
end
